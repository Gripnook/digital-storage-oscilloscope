package filter_parameters is

    constant HLP2_LENGTH : integer := 43;
    constant HLP2_PIPELINE_LENGTH : integer := 7;
    constant HLP4_LENGTH : integer := 86;
    constant HLP4_PIPELINE_LENGTH : integer := 8;
    constant HLP8_LENGTH : integer := 170;
    constant HLP8_PIPELINE_LENGTH : integer := 9;
    constant HLP16_LENGTH : integer := 339;
    constant HLP16_PIPELINE_LENGTH : integer := 10;

end package;
