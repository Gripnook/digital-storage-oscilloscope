package filter_parameters is
    
    constant HLP2_LENGTH : integer := 43;
    constant HLP4_LENGTH : integer := 86;
    constant HLP8_LENGTH : integer := 170;
    constant HLP16_LENGTH : integer := 339;

end package;
